module riscv #(parameter WIDTH=32)
(
);

endmodule