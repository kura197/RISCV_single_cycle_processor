`include "def.h";

module controller #() 
(
    input logic [`INSTR_BIT-1:0] kind,
    input logic [2:0] funct3,
    input logic [6:0] funct7
);
    
endmodule